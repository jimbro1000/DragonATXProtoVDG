`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:20:26 06/07/2025 
// Design Name: 
// Module Name:    RawSwitch 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RawSwitch(
    input [7:0] Data,
    input [3:0] Mode,
    input Css,
    input Clk,
    input Divider,
    input Load,    
    output [8:0] RGB
	 );



endmodule