module semi4Rom(
	input logic [7:0] inData,
	input logic [3:0] row,
	output logic [7:0] outData,
	output logic [3:0] colour
);

logic [7:0] semiData [0:3];

initial begin
	semiData[0] = 8'b11111111;
	semiData[1] = 8'b11110000;
	semiData[2] = 8'b00001111;
	semiData[3] = 8'b00000000;
end

logic [3:0] index;

always @(row, inData) begin
	case (row)
		0,1,2,3,4,5:
			index = inData[1:0];
		default:
			index = inData[3:2];
	endcase
	outData = semiData[index];
	colour = inData[6:4] + 1;
end

endmodule